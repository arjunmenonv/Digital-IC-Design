*** SPICE deck for cell INVERTER_LAYOUT{lay} from library EXPT1_2x
*** Created on Mon Sep 13, 2021 11:47:02
*** Last revised on Sat Sep 18, 2021 12:37:54
*** Written on Tue Sep 21, 2021 20:43:42 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: INVERTER_LAYOUT{lay}
Mnmos@1 OUT IN gnd gnd nmos L=0.022U W=0.088U AS=0.006P AD=0.009P PS=0.308U PD=0.396U
Mpmos@2 OUT IN vdd vdd pmos L=0.022U W=0.176U AS=0.012P AD=0.009P PS=0.484U PD=0.396U

* Spice Code nodes in cell cell 'INVERTER_LAYOUT{lay}'
.include "C:\Users\hp\OneDrive - smail.iitm.ac.in\Desktop\DIC\22nm_HP.pm"
v1 IN gnd pwl(0 0 10p 0 110p 0.8 1.1n 0.8 1.2n 0 2n 0)
v2 VDD gnd DC 0.8
.meas tran inv_fall_delay
+ trig v(in) val=0.4 cross=1
+ targ v(out) val=0.4 cross=1
.meas tran inv_rise_delay
+ trig v(in) val=0.4 cross=2
+ targ v(out) val=0.4 cross=2
.meas tran inv_trise
+ trig v(out) val=0.08 cross=2
+ targ v(out) val=0.72 cross=2
.meas tran inv_tfall
+ trig v(out) val=0.72 cross=1
+ targ v(out) val=0.08 cross=1
.tran 2.1n
.END
