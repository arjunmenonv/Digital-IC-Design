*** SPICE deck for cell NAND2_DELAY{sch} from library EXPT1_2x
*** Created on Sat Sep 18, 2021 21:01:20
*** Last revised on Wed Sep 22, 2021 17:40:28
*** Written on Wed Sep 22, 2021 17:41:09 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT EXPT1_2x__NAND2 FROM CELL NAND2{sch}
.SUBCKT EXPT1_2x__NAND2 A B gnd OUT vdd
Mnmos@0 OUT A net@6 gnd nmos L=0.022U W=0.176U
Mnmos@1 net@6 B gnd gnd nmos L=0.022U W=0.176U
Mpmos@0 vdd A OUT vdd pmos L=0.022U W=0.176U
Mpmos@1 vdd B OUT vdd pmos L=0.022U W=0.176U
.ENDS EXPT1_2x__NAND2

.global gnd vdd

*** TOP LEVEL CELL: NAND2_DELAY{sch}
XNAND2@12 vdd IN gnd OUT_PRIMARY vdd EXPT1_2x__NAND2
XNAND2@13 OUT_PRIMARY NAND2@13_B gnd NAND2@13_OUT vdd EXPT1_2x__NAND2
XNAND2@14 OUT_PRIMARY NAND2@14_B gnd NAND2@14_OUT vdd EXPT1_2x__NAND2
XNAND2@15 OUT_PRIMARY NAND2@15_B gnd NAND2@15_OUT vdd EXPT1_2x__NAND2
XNAND2@16 OUT_PRIMARY NAND2@16_B gnd NAND2@16_OUT vdd EXPT1_2x__NAND2
XNAND2@17 OUT_PRIMARY NAND2@17_B gnd NAND2@17_OUT vdd EXPT1_2x__NAND2
XNAND2@18 OUT_PRIMARY NAND2@18_B gnd NAND2@18_OUT vdd EXPT1_2x__NAND2
XNAND2@19 OUT_PRIMARY NAND2@19_B gnd NAND2@19_OUT vdd EXPT1_2x__NAND2
XNAND2@20 OUT_PRIMARY NAND2@20_B gnd NAND2@20_OUT vdd EXPT1_2x__NAND2

* Spice Code nodes in cell cell 'NAND2_DELAY{sch}'
*.include "C:\Users\hp\OneDrive - smail.iitm.ac.in\Desktop\DIC\22nm_HP.pm"
.include "/home/arjunmenonv/Arjun_acads/Year4/DigIC/22nm_HP.pm"
v1 IN gnd pwl(0 0 30p 0 130p 0.8 1.3n 0.8 1.4n 0 2n 0)
v2 VDD gnd DC 0.8
.meas tran inv_fall_delay
+ trig v(in) val=0.4 cross=1
+ targ v(out_primary) val=0.4 cross=1
.meas tran inv_rise_delay
+ trig v(in) val=0.4 cross=2
+ targ v(out_primary) val=0.4 cross=2
.meas tran inv_trise
+ trig v(out_primary) val=0.08 cross=2
+ targ v(out_primary) val=0.72 cross=2
.meas tran inv_tfall
+ trig v(out_primary) val=0.72 cross=1
+ targ v(out_primary) val=0.08 cross=1
.tran 2.1n
.END
