*** SPICE deck for cell FanOut_NAND2_1x{sch} from library Assign1
*** Created on Thu Sep 16, 2021 18:57:15
*** Last revised on Sun Sep 19, 2021 13:57:33
*** Written on Tue Sep 21, 2021 14:55:52 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Assign1__NAND2_1x FROM CELL NAND2_1x{sch}
.SUBCKT Assign1__NAND2_1x A B OUT
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT A net@14 gnd nmos L=0.022U W=0.088U
Mnmos@1 net@14 B gnd gnd nmos L=0.022U W=0.088U
Mpmos@0 vdd A OUT vdd pmos L=0.022U W=0.088U
Mpmos@1 vdd B OUT vdd pmos L=0.022U W=0.088U
.ENDS Assign1__NAND2_1x

.global gnd vdd

*** TOP LEVEL CELL: FanOut_NAND2_1x{sch}
XNAND2_1x@9 inp_a inp_b out Assign1__NAND2_1x
XNAND2_1x@10 NAND2_1x@10_A NAND2_1x@10_B net@92 Assign1__NAND2_1x
XNAND2_1x@11 NAND2_1x@11_A NAND2_1x@11_B net@93 Assign1__NAND2_1x
XNAND2_1x@12 NAND2_1x@12_A NAND2_1x@12_B net@94 Assign1__NAND2_1x
XNAND2_1x@13 NAND2_1x@13_A NAND2_1x@13_B net@95 Assign1__NAND2_1x
XNAND2_1x@14 NAND2_1x@14_A NAND2_1x@14_B net@96 Assign1__NAND2_1x
XNAND2_1x@15 NAND2_1x@15_A NAND2_1x@15_B net@97 Assign1__NAND2_1x
XNAND2_1x@16 NAND2_1x@16_A NAND2_1x@16_B net@98 Assign1__NAND2_1x
XNAND2_1x@17 NAND2_1x@17_A NAND2_1x@17_B net@99 Assign1__NAND2_1x

* Spice Code nodes in cell cell 'FanOut_NAND2_1x{sch}'
*.include "C:\Users\arjun\Desktop\DigIC\22nm_HP.pm"
.include "/home/arjunmenonv/Arjun_acads/Year4/DigIC/22nm_HP.pm"

.param vdd_voltage= 0.8
v1 vdd gnd {vdd_voltage}
v2 inp_a gnd PULSE(0 {vdd_voltage} 1n 100p 100p 400p 1n 3)
*v2 inp_a gnd {vdd_voltage}
*Period = 1n
*v3 inp_b gnd PULSE(0 {vdd_voltage} 1n 100p 100p 900p 2n 3)
v3 inp_b gnd {vdd_voltage}
*Period = 2n
.meas tran Trise
+trig v(out) val={0.1*vdd_voltage} cross=2
+targ v(out) val={0.9*vdd_voltage} cross=2
.meas tran Tfall
+trig v(out) val={0.9*vdd_voltage} cross=1
+targ v(out) val={0.1*vdd_voltage} cross=1
.meas tran rise_Delay
*+trig v(inp_b) val={0.5*vdd_voltage} cross=2
+trig v(inp_a) val={0.5*vdd_voltage} cross=2
+targ v(out) val={0.5*vdd_voltage} cross=2
.meas tran fall_Delay
*+trig v(inp_b) val={0.5*vdd_voltage} cross=1
+trig v(inp_a) val={0.5*vdd_voltage} cross=1
+targ v(out) val={0.5*vdd_voltage} cross=1
.tran 4.3n
.end
.END
