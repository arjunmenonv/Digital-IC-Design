*** SPICE deck for cell DUT_AND2_1x{sch} from library Assign1
*** Created on Thu Sep 16, 2021 21:59:11
*** Last revised on Tue Sep 21, 2021 14:54:03
*** Written on Tue Sep 21, 2021 14:54:09 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Assign1__INV_1x FROM CELL INV_1x{sch}
.SUBCKT Assign1__INV_1x INP OUT
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT INP gnd gnd nmos L=0.022U W=0.044U
Mpmos@0 vdd INP OUT vdd pmos L=0.022U W=0.088U
.ENDS Assign1__INV_1x

*** SUBCIRCUIT Assign1__NAND2_1x FROM CELL NAND2_1x{sch}
.SUBCKT Assign1__NAND2_1x A B OUT
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT A net@14 gnd nmos L=0.022U W=0.088U
Mnmos@1 net@14 B gnd gnd nmos L=0.022U W=0.088U
Mpmos@0 vdd A OUT vdd pmos L=0.022U W=0.088U
Mpmos@1 vdd B OUT vdd pmos L=0.022U W=0.088U
.ENDS Assign1__NAND2_1x

*** SUBCIRCUIT Assign1__AND2_1x FROM CELL AND2_1x{sch}
.SUBCKT Assign1__AND2_1x A B OUT Y
** GLOBAL gnd
** GLOBAL vdd
XINV_1x@1 Y OUT Assign1__INV_1x
XNAND2_1x@0 A B Y Assign1__NAND2_1x
.ENDS Assign1__AND2_1x

.global gnd vdd

*** TOP LEVEL CELL: DUT_AND2_1x{sch}
XAND2_1x@0 INP_A INP_B OUT AND2_1x@0_Y Assign1__AND2_1x

* Spice Code nodes in cell cell 'DUT_AND2_1x{sch}'
.include "/home/arjunmenonv/Arjun_acads/Year4/DigIC/22nm_HP.pm"
.param vdd_voltage= 0.8
v1 vdd gnd {vdd_voltage}
v2 inp_a gnd PULSE(0 {vdd_voltage} 1n 100p 100p 400p 1n 3) 
*Period = 1n
v3 inp_b gnd PULSE(0 {vdd_voltage} 1n 100p 100p 900p 2n 3) 
*Period = 2n
.tran 4.3n
.end
.END
